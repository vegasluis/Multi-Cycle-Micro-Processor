module pcplus(input[5:0] d,
output [5:0] q);

assign q = d + 6'd1; 

endmodule